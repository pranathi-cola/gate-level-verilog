module neo_matrix(input choice2, choice1, choice0, a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115, output outa0, outa1, outa2, outa3, outa4, outa5, outa6, outa7, outa8, outa9, outa10, outa11, outa12, outa13, outa14, outa15, outb0, outb1, outb2, outb3, outb4, outb5, outb6, outb7, outb8, outb9, outb10, outb11, outb12, outb13, outb14, outb15, outc0, outc1, outc2, outc3, outc4, outc5, outc6, outc7, outc8, outc9, outc10, outc11, outc12, outc13, outc14, outc15, outd0, outd1, outd2, outd3, outd4, outd5, outd6, outd7, outd8, outd9, outd10, outd11, outd12, outd13, outd14, outd15, oute0, oute1, oute2, oute3, oute4, oute5, oute6, oute7, oute8, oute9, oute10, oute11, oute12, oute13, oute14, oute15, outf0, outf1, outf2, outf3, outf4, outf5, outf6, outf7, outf8, outf9, outf10, outf11, outf12, outf13, outf14, outf15, outg0, outg1, outg2, outg3, outg4, outg5, outg6, outg7, outg8, outg9, outg10, outg11, outg12, outg13, outg14, outg15, outh0, outh1, outh2, outh3, outh4, outh5, outh6, outh7, outh8, outh9, outh10, outh11, outh12, outh13, outh14, outh15, outi0, outi1, outi2, outi3, outi4, outi5, outi6, outi7, outi8, outi9, outi10, outi11, outi12, outi13, outi14, outi15);

input choice2, choice1, choice0, a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115;
output outa0, outa1, outa2, outa3, outa4, outa5, outa6, outa7, outa8, outa9, outa10, outa11, outa12, outa13, outa14, outa15, outb0, outb1, outb2, outb3, outb4, outb5, outb6, outb7, outb8, outb9, outb10, outb11, outb12, outb13, outb14, outb15, outc0, outc1, outc2, outc3, outc4, outc5, outc6, outc7, outc8, outc9, outc10, outc11, outc12, outc13, outc14, outc15, outd0, outd1, outd2, outd3, outd4, outd5, outd6, outd7, outd8, outd9, outd10, outd11, outd12, outd13, outd14, outd15, oute0, oute1, oute2, oute3, oute4, oute5, oute6, oute7, oute8, oute9, oute10, oute11, oute12, oute13, oute14, oute15, outf0, outf1, outf2, outf3, outf4, outf5, outf6, outf7, outf8, outf9, outf10, outf11, outf12, outf13, outf14, outf15, outg0, outg1, outg2, outg3, outg4, outg5, outg6, outg7, outg8, outg9, outg10, outg11, outg12, outg13, outg14, outg15, outh0, outh1, outh2, outh3, outh4, outh5, outh6, outh7, outh8, outh9, outh10, outh11, outh12, outh13, outh14, outh15, outi0, outi1, outi2, outi3, outi4, outi5, outi6, outi7, outi8, outi9, outi10, outi11, outi12, outi13, outi14, outi15;
wire adda0, adda1, adda2, adda3, adda4, adda5, adda6, adda7, adda8, adda9, adda10, adda11, adda12, adda13, adda14, adda15, addb0, addb1, addb2, addb3, addb4, addb5, addb6, addb7, addb8, addb9, addb10, addb11, addb12, addb13, addb14, addb15, addc0, addc1, addc2, addc3, addc4, addc5, addc6, addc7, addc8, addc9, addc10, addc11, addc12, addc13, addc14, addc15, addd0, addd1, addd2, addd3, addd4, addd5, addd6, addd7, addd8, addd9, addd10, addd11, addd12, addd13, addd14, addd15, adde0, adde1, adde2, adde3, adde4, adde5, adde6, adde7, adde8, adde9, adde10, adde11, adde12, adde13, adde14, adde15, addf0, addf1, addf2, addf3, addf4, addf5, addf6, addf7, addf8, addf9, addf10, addf11, addf12, addf13, addf14, addf15, addg0, addg1, addg2, addg3, addg4, addg5, addg6, addg7, addg8, addg9, addg10, addg11, addg12, addg13, addg14, addg15, addh0, addh1, addh2, addh3, addh4, addh5, addh6, addh7, addh8, addh9, addh10, addh11, addh12, addh13, addh14, addh15, addi0, addi1, addi2, addi3, addi4, addi5, addi6, addi7, addi8, addi9, addi10, addi11, addi12, addi13, addi14, addi15;
wire suba0, suba1, suba2, suba3, suba4, suba5, suba6, suba7, suba8, suba9, suba10, suba11, suba12, suba13, suba14, suba15, subb0, subb1, subb2, subb3, subb4, subb5, subb6, subb7, subb8, subb9, subb10, subb11, subb12, subb13, subb14, subb15, subc0, subc1, subc2, subc3, subc4, subc5, subc6, subc7, subc8, subc9, subc10, subc11, subc12, subc13, subc14, subc15, subd0, subd1, subd2, subd3, subd4, subd5, subd6, subd7, subd8, subd9, subd10, subd11, subd12, subd13, subd14, subd15, sube0, sube1, sube2, sube3, sube4, sube5, sube6, sube7, sube8, sube9, sube10, sube11, sube12, sube13, sube14, sube15, subf0, subf1, subf2, subf3, subf4, subf5, subf6, subf7, subf8, subf9, subf10, subf11, subf12, subf13, subf14, subf15, subg0, subg1, subg2, subg3, subg4, subg5, subg6, subg7, subg8, subg9, subg10, subg11, subg12, subg13, subg14, subg15, subh0, subh1, subh2, subh3, subh4, subh5, subh6, subh7, subh8, subh9, subh10, subh11, subh12, subh13, subh14, subh15, subi0, subi1, subi2, subi3, subi4, subi5, subi6, subi7, subi8, subi9, subi10, subi11, subi12, subi13, subi14, subi15;
wire multia0, multia1, multia2, multia3, multia4, multia5, multia6, multia7, multia8, multia9, multia10, multia11, multia12, multia13, multia14, multia15, multib0, multib1, multib2, multib3, multib4, multib5, multib6, multib7, multib8, multib9, multib10, multib11, multib12, multib13, multib14, multib15, multic0, multic1, multic2, multic3, multic4, multic5, multic6, multic7, multic8, multic9, multic10, multic11, multic12, multic13, multic14, multic15, multid0, multid1, multid2, multid3, multid4, multid5, multid6, multid7, multid8, multid9, multid10, multid11, multid12, multid13, multid14, multid15, multie0, multie1, multie2, multie3, multie4, multie5, multie6, multie7, multie8, multie9, multie10, multie11, multie12, multie13, multie14, multie15, multif0, multif1, multif2, multif3, multif4, multif5, multif6, multif7, multif8, multif9, multif10, multif11, multif12, multif13, multif14, multif15, multig0, multig1, multig2, multig3, multig4, multig5, multig6, multig7, multig8, multig9, multig10, multig11, multig12, multig13, multig14, multig15, multih0, multih1, multih2, multih3, multih4, multih5, multih6, multih7, multih8, multih9, multih10, multih11, multih12, multih13, multih14, multih15, multii0, multii1, multii2, multii3, multii4, multii5, multii6, multii7, multii8, multii9, multii10, multii11, multii12, multii13, multii14, multii15;
wire diva0, diva1, diva2, diva3, diva4, diva5, diva6, diva7, diva8, diva9, diva10, diva11, diva12, diva13, diva14, diva15, divb0, divb1, divb2, divb3, divb4, divb5, divb6, divb7, divb8, divb9, divb10, divb11, divb12, divb13, divb14, divb15, divc0, divc1, divc2, divc3, divc4, divc5, divc6, divc7, divc8, divc9, divc10, divc11, divc12, divc13, divc14, divc15, divd0, divd1, divd2, divd3, divd4, divd5, divd6, divd7, divd8, divd9, divd10, divd11, divd12, divd13, divd14, divd15, dive0, dive1, dive2, dive3, dive4, dive5, dive6, dive7, dive8, dive9, dive10, dive11, dive12, dive13, dive14, dive15, divf0, divf1, divf2, divf3, divf4, divf5, divf6, divf7, divf8, divf9, divf10, divf11, divf12, divf13, divf14, divf15, divg0, divg1, divg2, divg3, divg4, divg5, divg6, divg7, divg8, divg9, divg10, divg11, divg12, divg13, divg14, divg15, divh0, divh1, divh2, divh3, divh4, divh5, divh6, divh7, divh8, divh9, divh10, divh11, divh12, divh13, divh14, divh15, divi0, divi1, divi2, divi3, divi4, divi5, divi6, divi7, divi8, divi9, divi10, divi11, divi12, divi13, divi14, divi15;
wire inva0, inva1, inva2, inva3, inva4, inva5, inva6, inva7, inva8, inva9, inva10, inva11, inva12, inva13, inva14, inva15, invb0, invb1, invb2, invb3, invb4, invb5, invb6, invb7, invb8, invb9, invb10, invb11, invb12, invb13, invb14, invb15, invc0, invc1, invc2, invc3, invc4, invc5, invc6, invc7, invc8, invc9, invc10, invc11, invc12, invc13, invc14, invc15, invd0, invd1, invd2, invd3, invd4, invd5, invd6, invd7, invd8, invd9, invd10, invd11, invd12, invd13, invd14, invd15, inve0, inve1, inve2, inve3, inve4, inve5, inve6, inve7, inve8, inve9, inve10, inve11, inve12, inve13, inve14, inve15, invf0, invf1, invf2, invf3, invf4, invf5, invf6, invf7, invf8, invf9, invf10, invf11, invf12, invf13, invf14, invf15, invg0, invg1, invg2, invg3, invg4, invg5, invg6, invg7, invg8, invg9, invg10, invg11, invg12, invg13, invg14, invg15, invh0, invh1, invh2, invh3, invh4, invh5, invh6, invh7, invh8, invh9, invh10, invh11, invh12, invh13, invh14, invh15, invi0, invi1, invi2, invi3, invi4, invi5, invi6, invi7, invi8, invi9, invi10, invi11, invi12, invi13, invi14, invi15;

matrix_adder matrix1(a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115, adda0, adda1, adda2, adda3, adda4, adda5, adda6, adda7, adda8, adda9, adda10, adda11, adda12, adda13, adda14, adda15, addb0, addb1, addb2, addb3, addb4, addb5, addb6, addb7, addb8, addb9, addb10, addb11, addb12, addb13, addb14, addb15, addc0, addc1, addc2, addc3, addc4, addc5, addc6, addc7, addc8, addc9, addc10, addc11, addc12, addc13, addc14, addc15, addd0, addd1, addd2, addd3, addd4, addd5, addd6, addd7, addd8, addd9, addd10, addd11, addd12, addd13, addd14, addd15, adde0, adde1, adde2, adde3, adde4, adde5, adde6, adde7, adde8, adde9, adde10, adde11, adde12, adde13, adde14, adde15, addf0, addf1, addf2, addf3, addf4, addf5, addf6, addf7, addf8, addf9, addf10, addf11, addf12, addf13, addf14, addf15, addg0, addg1, addg2, addg3, addg4, addg5, addg6, addg7, addg8, addg9, addg10, addg11, addg12, addg13, addg14, addg15, addh0, addh1, addh2, addh3, addh4, addh5, addh6, addh7, addh8, addh9, addh10, addh11, addh12, addh13, addh14, addh15, addi0, addi1, addi2, addi3, addi4, addi5, addi6, addi7, addi8, addi9, addi10, addi11, addi12, addi13, addi14, addi15);
matrix_subtractor matrix2(a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115, suba0, suba1, suba2, suba3, suba4, suba5, suba6, suba7, suba8, suba9, suba10, suba11, suba12, suba13, suba14, suba15, subb0, subb1, subb2, subb3, subb4, subb5, subb6, subb7, subb8, subb9, subb10, subb11, subb12, subb13, subb14, subb15, subc0, subc1, subc2, subc3, subc4, subc5, subc6, subc7, subc8, subc9, subc10, subc11, subc12, subc13, subc14, subc15, subd0, subd1, subd2, subd3, subd4, subd5, subd6, subd7, subd8, subd9, subd10, subd11, subd12, subd13, subd14, subd15, sube0, sube1, sube2, sube3, sube4, sube5, sube6, sube7, sube8, sube9, sube10, sube11, sube12, sube13, sube14, sube15, subf0, subf1, subf2, subf3, subf4, subf5, subf6, subf7, subf8, subf9, subf10, subf11, subf12, subf13, subf14, subf15, subg0, subg1, subg2, subg3, subg4, subg5, subg6, subg7, subg8, subg9, subg10, subg11, subg12, subg13, subg14, subg15, subh0, subh1, subh2, subh3, subh4, subh5, subh6, subh7, subh8, subh9, subh10, subh11, subh12, subh13, subh14, subh15, subi0, subi1, subi2, subi3, subi4, subi5, subi6, subi7, subi8, subi9, subi10, subi11, subi12, subi13, subi14, subi15);
matrix_multiply matrix3(a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115, multia0, multia1, multia2, multia3, multia4, multia5, multia6, multia7, multia8, multia9, multia10, multia11, multia12, multia13, multia14, multia15, multib0, multib1, multib2, multib3, multib4, multib5, multib6, multib7, multib8, multib9, multib10, multib11, multib12, multib13, multib14, multib15, multic0, multic1, multic2, multic3, multic4, multic5, multic6, multic7, multic8, multic9, multic10, multic11, multic12, multic13, multic14, multic15, multid0, multid1, multid2, multid3, multid4, multid5, multid6, multid7, multid8, multid9, multid10, multid11, multid12, multid13, multid14, multid15, multie0, multie1, multie2, multie3, multie4, multie5, multie6, multie7, multie8, multie9, multie10, multie11, multie12, multie13, multie14, multie15, multif0, multif1, multif2, multif3, multif4, multif5, multif6, multif7, multif8, multif9, multif10, multif11, multif12, multif13, multif14, multif15, multig0, multig1, multig2, multig3, multig4, multig5, multig6, multig7, multig8, multig9, multig10, multig11, multig12, multig13, multig14, multig15, multih0, multih1, multih2, multih3, multih4, multih5, multih6, multih7, multih8, multih9, multih10, multih11, multih12, multih13, multih14, multih15, multii0, multii1, multii2, multii3, multii4, multii5, multii6, multii7, multii8, multii9, multii10, multii11, multii12, multii13, multii14, multii15);
matrix_scalar_division matrix4(a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115, diva0, diva1, diva2, diva3, diva4, diva5, diva6, diva7, diva8, diva9, diva10, diva11, diva12, diva13, diva14, diva15, divb0, divb1, divb2, divb3, divb4, divb5, divb6, divb7, divb8, divb9, divb10, divb11, divb12, divb13, divb14, divb15, divc0, divc1, divc2, divc3, divc4, divc5, divc6, divc7, divc8, divc9, divc10, divc11, divc12, divc13, divc14, divc15, divd0, divd1, divd2, divd3, divd4, divd5, divd6, divd7, divd8, divd9, divd10, divd11, divd12, divd13, divd14, divd15, dive0, dive1, dive2, dive3, dive4, dive5, dive6, dive7, dive8, dive9, dive10, dive11, dive12, dive13, dive14, dive15, divf0, divf1, divf2, divf3, divf4, divf5, divf6, divf7, divf8, divf9, divf10, divf11, divf12, divf13, divf14, divf15, divg0, divg1, divg2, divg3, divg4, divg5, divg6, divg7, divg8, divg9, divg10, divg11, divg12, divg13, divg14, divg15, divh0, divh1, divh2, divh3, divh4, divh5, divh6, divh7, divh8, divh9, divh10, divh11, divh12, divh13, divh14, divh15, divi0, divi1, divi2, divi3, divi4, divi5, divi6, divi7, divi8, divi9, divi10, divi11, divi12, divi13, divi14, divi15);
matrix_division matrix5(a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115, inva0, inva1, inva2, inva3, inva4, inva5, inva6, inva7, inva8, inva9, inva10, inva11, inva12, inva13, inva14, inva15, invb0, invb1, invb2, invb3, invb4, invb5, invb6, invb7, invb8, invb9, invb10, invb11, invb12, invb13, invb14, invb15, invc0, invc1, invc2, invc3, invc4, invc5, invc6, invc7, invc8, invc9, invc10, invc11, invc12, invc13, invc14, invc15, invd0, invd1, invd2, invd3, invd4, invd5, invd6, invd7, invd8, invd9, invd10, invd11, invd12, invd13, invd14, invd15, inve0, inve1, inve2, inve3, inve4, inve5, inve6, inve7, inve8, inve9, inve10, inve11, inve12, inve13, inve14, inve15, invf0, invf1, invf2, invf3, invf4, invf5, invf6, invf7, invf8, invf9, invf10, invf11, invf12, invf13, invf14, invf15, invg0, invg1, invg2, invg3, invg4, invg5, invg6, invg7, invg8, invg9, invg10, invg11, invg12, invg13, invg14, invg15, invh0, invh1, invh2, invh3, invh4, invh5, invh6, invh7, invh8, invh9, invh10, invh11, invh12, invh13, invh14, invh15, invi0, invi1, invi2, invi3, invi4, invi5, invi6, invi7, invi8, invi9, invi10, invi11, invi12, invi13, invi14, invi15);

lol1 l00(choice2, choice1, choice0, adda0, suba0, multia0, diva0, inva0, outa0);
lol1 l01(choice2, choice1, choice0, adda1, suba1, multia1, diva1, inva1, outa1);
lol1 l02(choice2, choice1, choice0, adda2, suba2, multia2, diva2, inva2, outa2);
lol1 l03(choice2, choice1, choice0, adda3, suba3, multia3, diva3, inva3, outa3);
lol1 l04(choice2, choice1, choice0, adda4, suba4, multia4, diva4, inva4, outa4);
lol1 l05(choice2, choice1, choice0, adda5, suba5, multia5, diva5, inva5, outa5);
lol1 l06(choice2, choice1, choice0, adda6, suba6, multia6, diva6, inva6, outa6);
lol1 l07(choice2, choice1, choice0, adda7, suba7, multia7, diva7, inva7, outa7);
lol1 l08(choice2, choice1, choice0, adda8, suba8, multia8, diva8, inva8, outa8);
lol1 l09(choice2, choice1, choice0, adda9, suba9, multia9, diva9, inva9, outa9);
lol1 l010(choice2, choice1, choice0, adda10, suba10, multia10, diva10, inva10, outa10);
lol1 l011(choice2, choice1, choice0, adda11, suba11, multia11, diva11, inva11, outa11);
lol1 l012(choice2, choice1, choice0, adda12, suba12, multia12, diva12, inva12, outa12);
lol1 l013(choice2, choice1, choice0, adda13, suba13, multia13, diva13, inva13, outa13);
lol1 l014(choice2, choice1, choice0, adda14, suba14, multia14, diva14, inva14, outa14);
lol1 l015(choice2, choice1, choice0, adda15, suba15, multia15, diva15, inva15, outa15);

lol1 l10(choice2, choice1, choice0, addb0, subb0, multib0, divb0, invb0, outb0);
lol1 l11(choice2, choice1, choice0, addb1, subb1, multib1, divb1, invb1, outb1);
lol1 l12(choice2, choice1, choice0, addb2, subb2, multib2, divb2, invb2, outb2);
lol1 l13(choice2, choice1, choice0, addb3, subb3, multib3, divb3, invb3, outb3);
lol1 l14(choice2, choice1, choice0, addb4, subb4, multib4, divb4, invb4, outb4);
lol1 l15(choice2, choice1, choice0, addb5, subb5, multib5, divb5, invb5, outb5);
lol1 l16(choice2, choice1, choice0, addb6, subb6, multib6, divb6, invb6, outb6);
lol1 l17(choice2, choice1, choice0, addb7, subb7, multib7, divb7, invb7, outb7);
lol1 l18(choice2, choice1, choice0, addb8, subb8, multib8, divb8, invb8, outb8);
lol1 l19(choice2, choice1, choice0, addb9, subb9, multib9, divb9, invb9, outb9);
lol1 l110(choice2, choice1, choice0, addb10, subb10, multib10, divb10, invb10, outb10);
lol1 l111(choice2, choice1, choice0, addb11, subb11, multib11, divb11, invb11, outb11);
lol1 l112(choice2, choice1, choice0, addb12, subb12, multib12, divb12, invb12, outb12);
lol1 l113(choice2, choice1, choice0, addb13, subb13, multib13, divb13, invb13, outb13);
lol1 l114(choice2, choice1, choice0, addb14, subb14, multib14, divb14, invb14, outb14);
lol1 l115(choice2, choice1, choice0, addb15, subb15, multib15, divb15, invb15, outb15);

lol1 l20(choice2, choice1, choice0, addc0, subc0, multic0, divc0, invc0, outc0);
lol1 l21(choice2, choice1, choice0, addc1, subc1, multic1, divc1, invc1, outc1);
lol1 l22(choice2, choice1, choice0, addc2, subc2, multic2, divc2, invc2, outc2);
lol1 l23(choice2, choice1, choice0, addc3, subc3, multic3, divc3, invc3, outc3);
lol1 l24(choice2, choice1, choice0, addc4, subc4, multic4, divc4, invc4, outc4);
lol1 l25(choice2, choice1, choice0, addc5, subc5, multic5, divc5, invc5, outc5);
lol1 l26(choice2, choice1, choice0, addc6, subc6, multic6, divc6, invc6, outc6);
lol1 l27(choice2, choice1, choice0, addc7, subc7, multic7, divc7, invc7, outc7);
lol1 l28(choice2, choice1, choice0, addc8, subc8, multic8, divc8, invc8, outc8);
lol1 l29(choice2, choice1, choice0, addc9, subc9, multic9, divc9, invc9, outc9);
lol1 l210(choice2, choice1, choice0, addc10, subc10, multic10, divc10, invc10, outc10);
lol1 l211(choice2, choice1, choice0, addc11, subc11, multic11, divc11, invc11, outc11);
lol1 l212(choice2, choice1, choice0, addc12, subc12, multic12, divc12, invc12, outc12);
lol1 l213(choice2, choice1, choice0, addc13, subc13, multic13, divc13, invc13, outc13);
lol1 l214(choice2, choice1, choice0, addc14, subc14, multic14, divc14, invc14, outc14);
lol1 l215(choice2, choice1, choice0, addc15, subc15, multic15, divc15, invc15, outc15);

lol1 l30(choice2, choice1, choice0, addd0, subd0, multid0, divd0, invd0, outd0);
lol1 l31(choice2, choice1, choice0, addd1, subd1, multid1, divd1, invd1, outd1);
lol1 l32(choice2, choice1, choice0, addd2, subd2, multid2, divd2, invd2, outd2);
lol1 l33(choice2, choice1, choice0, addd3, subd3, multid3, divd3, invd3, outd3);
lol1 l34(choice2, choice1, choice0, addd4, subd4, multid4, divd4, invd4, outd4);
lol1 l35(choice2, choice1, choice0, addd5, subd5, multid5, divd5, invd5, outd5);
lol1 l36(choice2, choice1, choice0, addd6, subd6, multid6, divd6, invd6, outd6);
lol1 l37(choice2, choice1, choice0, addd7, subd7, multid7, divd7, invd7, outd7);
lol1 l38(choice2, choice1, choice0, addd8, subd8, multid8, divd8, invd8, outd8);
lol1 l39(choice2, choice1, choice0, addd9, subd9, multid9, divd9, invd9, outd9);
lol1 l310(choice2, choice1, choice0, addd10, subd10, multid10, divd10, invd10, outd10);
lol1 l311(choice2, choice1, choice0, addd11, subd11, multid11, divd11, invd11, outd11);
lol1 l312(choice2, choice1, choice0, addd12, subd12, multid12, divd12, invd12, outd12);
lol1 l313(choice2, choice1, choice0, addd13, subd13, multid13, divd13, invd13, outd13);
lol1 l314(choice2, choice1, choice0, addd14, subd14, multid14, divd14, invd14, outd14);
lol1 l315(choice2, choice1, choice0, addd15, subd15, multid15, divd15, invd15, outd15);

lol1 l40(choice2, choice1, choice0, adde0, sube0, multie0, dive0, inve0, oute0);
lol1 l41(choice2, choice1, choice0, adde1, sube1, multie1, dive1, inve1, oute1);
lol1 l42(choice2, choice1, choice0, adde2, sube2, multie2, dive2, inve2, oute2);
lol1 l43(choice2, choice1, choice0, adde3, sube3, multie3, dive3, inve3, oute3);
lol1 l44(choice2, choice1, choice0, adde4, sube4, multie4, dive4, inve4, oute4);
lol1 l45(choice2, choice1, choice0, adde5, sube5, multie5, dive5, inve5, oute5);
lol1 l46(choice2, choice1, choice0, adde6, sube6, multie6, dive6, inve6, oute6);
lol1 l47(choice2, choice1, choice0, adde7, sube7, multie7, dive7, inve7, oute7);
lol1 l48(choice2, choice1, choice0, adde8, sube8, multie8, dive8, inve8, oute8);
lol1 l49(choice2, choice1, choice0, adde9, sube9, multie9, dive9, inve9, oute9);
lol1 l410(choice2, choice1, choice0, adde10, sube10, multie10, dive10, inve10, oute10);
lol1 l411(choice2, choice1, choice0, adde11, sube11, multie11, dive11, inve11, oute11);
lol1 l412(choice2, choice1, choice0, adde12, sube12, multie12, dive12, inve12, oute12);
lol1 l413(choice2, choice1, choice0, adde13, sube13, multie13, dive13, inve13, oute13);
lol1 l414(choice2, choice1, choice0, adde14, sube14, multie14, dive14, inve14, oute14);
lol1 l415(choice2, choice1, choice0, adde15, sube15, multie15, dive15, inve15, oute15);

lol1 l50(choice2, choice1, choice0, addf0, subf0, multif0, divf0, invf0, outf0);
lol1 l51(choice2, choice1, choice0, addf1, subf1, multif1, divf1, invf1, outf1);
lol1 l52(choice2, choice1, choice0, addf2, subf2, multif2, divf2, invf2, outf2);
lol1 l53(choice2, choice1, choice0, addf3, subf3, multif3, divf3, invf3, outf3);
lol1 l54(choice2, choice1, choice0, addf4, subf4, multif4, divf4, invf4, outf4);
lol1 l55(choice2, choice1, choice0, addf5, subf5, multif5, divf5, invf5, outf5);
lol1 l56(choice2, choice1, choice0, addf6, subf6, multif6, divf6, invf6, outf6);
lol1 l57(choice2, choice1, choice0, addf7, subf7, multif7, divf7, invf7, outf7);
lol1 l58(choice2, choice1, choice0, addf8, subf8, multif8, divf8, invf8, outf8);
lol1 l59(choice2, choice1, choice0, addf9, subf9, multif9, divf9, invf9, outf9);
lol1 l510(choice2, choice1, choice0, addf10, subf10, multif10, divf10, invf10, outf10);
lol1 l511(choice2, choice1, choice0, addf11, subf11, multif11, divf11, invf11, outf11);
lol1 l512(choice2, choice1, choice0, addf12, subf12, multif12, divf12, invf12, outf12);
lol1 l513(choice2, choice1, choice0, addf13, subf13, multif13, divf13, invf13, outf13);
lol1 l514(choice2, choice1, choice0, addf14, subf14, multif14, divf14, invf14, outf14);
lol1 l515(choice2, choice1, choice0, addf15, subf15, multif15, divf15, invf15, outf15);

lol1 l60(choice2, choice1, choice0, addg0, subg0, multig0, divg0, invg0, outg0);
lol1 l61(choice2, choice1, choice0, addg1, subg1, multig1, divg1, invg1, outg1);
lol1 l62(choice2, choice1, choice0, addg2, subg2, multig2, divg2, invg2, outg2);
lol1 l63(choice2, choice1, choice0, addg3, subg3, multig3, divg3, invg3, outg3);
lol1 l64(choice2, choice1, choice0, addg4, subg4, multig4, divg4, invg4, outg4);
lol1 l65(choice2, choice1, choice0, addg5, subg5, multig5, divg5, invg5, outg5);
lol1 l66(choice2, choice1, choice0, addg6, subg6, multig6, divg6, invg6, outg6);
lol1 l67(choice2, choice1, choice0, addg7, subg7, multig7, divg7, invg7, outg7);
lol1 l68(choice2, choice1, choice0, addg8, subg8, multig8, divg8, invg8, outg8);
lol1 l69(choice2, choice1, choice0, addg9, subg9, multig9, divg9, invg9, outg9);
lol1 l610(choice2, choice1, choice0, addg10, subg10, multig10, divg10, invg10, outg10);
lol1 l611(choice2, choice1, choice0, addg11, subg11, multig11, divg11, invg11, outg11);
lol1 l612(choice2, choice1, choice0, addg12, subg12, multig12, divg12, invg12, outg12);
lol1 l613(choice2, choice1, choice0, addg13, subg13, multig13, divg13, invg13, outg13);
lol1 l614(choice2, choice1, choice0, addg14, subg14, multig14, divg14, invg14, outg14);
lol1 l615(choice2, choice1, choice0, addg15, subg15, multig15, divg15, invg15, outg15);

lol1 l70(choice2, choice1, choice0, addh0, subh0, multih0, divh0, invh0, outh0);
lol1 l71(choice2, choice1, choice0, addh1, subh1, multih1, divh1, invh1, outh1);
lol1 l72(choice2, choice1, choice0, addh2, subh2, multih2, divh2, invh2, outh2);
lol1 l73(choice2, choice1, choice0, addh3, subh3, multih3, divh3, invh3, outh3);
lol1 l74(choice2, choice1, choice0, addh4, subh4, multih4, divh4, invh4, outh4);
lol1 l75(choice2, choice1, choice0, addh5, subh5, multih5, divh5, invh5, outh5);
lol1 l76(choice2, choice1, choice0, addh6, subh6, multih6, divh6, invh6, outh6);
lol1 l77(choice2, choice1, choice0, addh7, subh7, multih7, divh7, invh7, outh7);
lol1 l78(choice2, choice1, choice0, addh8, subh8, multih8, divh8, invh8, outh8);
lol1 l79(choice2, choice1, choice0, addh9, subh9, multih9, divh9, invh9, outh9);
lol1 l710(choice2, choice1, choice0, addh10, subh10, multih10, divh10, invh10, outh10);
lol1 l711(choice2, choice1, choice0, addh11, subh11, multih11, divh11, invh11, outh11);
lol1 l712(choice2, choice1, choice0, addh12, subh12, multih12, divh12, invh12, outh12);
lol1 l713(choice2, choice1, choice0, addh13, subh13, multih13, divh13, invh13, outh13);
lol1 l714(choice2, choice1, choice0, addh14, subh14, multih14, divh14, invh14, outh14);
lol1 l715(choice2, choice1, choice0, addh15, subh15, multih15, divh15, invh15, outh15);

lol1 l80(choice2, choice1, choice0, addi0, subi0, multii0, divi0, invi0, outi0);
lol1 l81(choice2, choice1, choice0, addi1, subi1, multii1, divi1, invi1, outi1);
lol1 l82(choice2, choice1, choice0, addi2, subi2, multii2, divi2, invi2, outi2);
lol1 l83(choice2, choice1, choice0, addi3, subi3, multii3, divi3, invi3, outi3);
lol1 l84(choice2, choice1, choice0, addi4, subi4, multii4, divi4, invi4, outi4);
lol1 l85(choice2, choice1, choice0, addi5, subi5, multii5, divi5, invi5, outi5);
lol1 l86(choice2, choice1, choice0, addi6, subi6, multii6, divi6, invi6, outi6);
lol1 l87(choice2, choice1, choice0, addi7, subi7, multii7, divi7, invi7, outi7);
lol1 l88(choice2, choice1, choice0, addi8, subi8, multii8, divi8, invi8, outi8);
lol1 l89(choice2, choice1, choice0, addi9, subi9, multii9, divi9, invi9, outi9);
lol1 l810(choice2, choice1, choice0, addi10, subi10, multii10, divi10, invi10, outi10);
lol1 l811(choice2, choice1, choice0, addi11, subi11, multii11, divi11, invi11, outi11);
lol1 l812(choice2, choice1, choice0, addi12, subi12, multii12, divi12, invi12, outi12);
lol1 l813(choice2, choice1, choice0, addi13, subi13, multii13, divi13, invi13, outi13);
lol1 l814(choice2, choice1, choice0, addi14, subi14, multii14, divi14, invi14, outi14);
lol1 l815(choice2, choice1, choice0, addi15, subi15, multii15, divi15, invi15, outi15);

endmodule
