module matrix_adder(input a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115, output outa0, outa1, outa2, outa3, outa4, outa5, outa6, outa7, outa8, outa9, outa10, outa11, outa12, outa13, outa14, outa15, outb0, outb1, outb2, outb3, outb4, outb5, outb6, outb7, outb8, outb9, outb10, outb11, outb12, outb13, outb14, outb15, outc0, outc1, outc2, outc3, outc4, outc5, outc6, outc7, outc8, outc9, outc10, outc11, outc12, outc13, outc14, outc15, outd0, outd1, outd2, outd3, outd4, outd5, outd6, outd7, outd8, outd9, outd10, outd11, outd12, outd13, outd14, outd15, oute0, oute1, oute2, oute3, oute4, oute5, oute6, oute7, oute8, oute9, oute10, oute11, oute12, oute13, oute14, oute15, outf0, outf1, outf2, outf3, outf4, outf5, outf6, outf7, outf8, outf9, outf10, outf11, outf12, outf13, outf14, outf15, outg0, outg1, outg2, outg3, outg4, outg5, outg6, outg7, outg8, outg9, outg10, outg11, outg12, outg13, outg14, outg15, outh0, outh1, outh2, outh3, outh4, outh5, outh6, outh7, outh8, outh9, outh10, outh11, outh12, outh13, outh14, outh15, outi0, outi1, outi2, outi3, outi4, outi5, outi6, outi7, outi8, outi9, outi10, outi11, outi12, outi13, outi14, outi15);

input a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115;
output outa0, outa1, outa2, outa3, outa4, outa5, outa6, outa7, outa8, outa9, outa10, outa11, outa12, outa13, outa14, outa15, outb0, outb1, outb2, outb3, outb4, outb5, outb6, outb7, outb8, outb9, outb10, outb11, outb12, outb13, outb14, outb15, outc0, outc1, outc2, outc3, outc4, outc5, outc6, outc7, outc8, outc9, outc10, outc11, outc12, outc13, outc14, outc15, outd0, outd1, outd2, outd3, outd4, outd5, outd6, outd7, outd8, outd9, outd10, outd11, outd12, outd13, outd14, outd15, oute0, oute1, oute2, oute3, oute4, oute5, oute6, oute7, oute8, oute9, oute10, oute11, oute12, oute13, oute14, oute15, outf0, outf1, outf2, outf3, outf4, outf5, outf6, outf7, outf8, outf9, outf10, outf11, outf12, outf13, outf14, outf15, outg0, outg1, outg2, outg3, outg4, outg5, outg6, outg7, outg8, outg9, outg10, outg11, outg12, outg13, outg14, outg15, outh0, outh1, outh2, outh3, outh4, outh5, outh6, outh7, outh8, outh9, outh10, outh11, outh12, outh13, outh14, outh15, outi0, outi1, outi2, outi3, outi4, outi5, outi6, outi7, outi8, outi9, outi10, outi11, outi12, outi13, outi14, outi15;

element_add element1(a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, outa0, outa1, outa2, outa3, outa4, outa5, outa6, outa7, outa8, outa9, outa10, outa11, outa12, outa13, outa14, outa15);
element_add element2(b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, outb0, outb1, outb2, outb3, outb4, outb5, outb6, outb7, outb8, outb9, outb10, outb11, outb12, outb13, outb14, outb15);
element_add element3(c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, outc0, outc1, outc2, outc3, outc4, outc5, outc6, outc7, outc8, outc9, outc10, outc11, outc12, outc13, outc14, outc15);
element_add element4(d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, outd0, outd1, outd2, outd3, outd4, outd5, outd6, outd7, outd8, outd9, outd10, outd11, outd12, outd13, outd14, outd15);
element_add element5(e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, oute0, oute1, oute2, oute3, oute4, oute5, oute6, oute7, oute8, oute9, oute10, oute11, oute12, oute13, oute14, oute15);
element_add element6(f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, outf0, outf1, outf2, outf3, outf4, outf5, outf6, outf7, outf8, outf9, outf10, outf11, outf12, outf13, outf14, outf15);
element_add element7(g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, outg0, outg1, outg2, outg3, outg4, outg5, outg6, outg7, outg8, outg9, outg10, outg11, outg12, outg13, outg14, outg15);
element_add element8(h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, outh0, outh1, outh2, outh3, outh4, outh5, outh6, outh7, outh8, outh9, outh10, outh11, outh12, outh13, outh14, outh15);
element_add element9(i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115, outi0, outi1, outi2, outi3, outi4, outi5, outi6, outi7, outi8, outi9, outi10, outi11, outi12, outi13, outi14, outi15);

endmodule
