module matrix_division(input a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115, output outa0, outa1, outa2, outa3, outa4, outa5, outa6, outa7, outa8, outa9, outa10, outa11, outa12, outa13, outa14, outa15, outb0, outb1, outb2, outb3, outb4, outb5, outb6, outb7, outb8, outb9, outb10, outb11, outb12, outb13, outb14, outb15, outc0, outc1, outc2, outc3, outc4, outc5, outc6, outc7, outc8, outc9, outc10, outc11, outc12, outc13, outc14, outc15, outd0, outd1, outd2, outd3, outd4, outd5, outd6, outd7, outd8, outd9, outd10, outd11, outd12, outd13, outd14, outd15, oute0, oute1, oute2, oute3, oute4, oute5, oute6, oute7, oute8, oute9, oute10, oute11, oute12, oute13, oute14, oute15, outf0, outf1, outf2, outf3, outf4, outf5, outf6, outf7, outf8, outf9, outf10, outf11, outf12, outf13, outf14, outf15, outg0, outg1, outg2, outg3, outg4, outg5, outg6, outg7, outg8, outg9, outg10, outg11, outg12, outg13, outg14, outg15, outh0, outh1, outh2, outh3, outh4, outh5, outh6, outh7, outh8, outh9, outh10, outh11, outh12, outh13, outh14, outh15, outi0, outi1, outi2, outi3, outi4, outi5, outi6, outi7, outi8, outi9, outi10, outi11, outi12, outi13, outi14, outi15);

input a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115;
output outa0, outa1, outa2, outa3, outa4, outa5, outa6, outa7, outa8, outa9, outa10, outa11, outa12, outa13, outa14, outa15, outb0, outb1, outb2, outb3, outb4, outb5, outb6, outb7, outb8, outb9, outb10, outb11, outb12, outb13, outb14, outb15, outc0, outc1, outc2, outc3, outc4, outc5, outc6, outc7, outc8, outc9, outc10, outc11, outc12, outc13, outc14, outc15, outd0, outd1, outd2, outd3, outd4, outd5, outd6, outd7, outd8, outd9, outd10, outd11, outd12, outd13, outd14, outd15, oute0, oute1, oute2, oute3, oute4, oute5, oute6, oute7, oute8, oute9, oute10, oute11, oute12, oute13, oute14, oute15, outf0, outf1, outf2, outf3, outf4, outf5, outf6, outf7, outf8, outf9, outf10, outf11, outf12, outf13, outf14, outf15, outg0, outg1, outg2, outg3, outg4, outg5, outg6, outg7, outg8, outg9, outg10, outg11, outg12, outg13, outg14, outg15, outh0, outh1, outh2, outh3, outh4, outh5, outh6, outh7, outh8, outh9, outh10, outh11, outh12, outh13, outh14, outh15, outi0, outi1, outi2, outi3, outi4, outi5, outi6, outi7, outi8, outi9, outi10, outi11, outi12, outi13, outi14, outi15;
wire a20, a21, a22, a23, b20, b21, b22, b23, c20, c21, c22, c23, d20, d21, d22, d23, e20, e21, e22, e23, f20, f21, f22, f23, g20, g21, g22, g23, h20, h21, h22, h23, i20, i21, i22, i23, a30, a31, a32, a33, b30, b31, b32, b33, c30, c31, c32, c33, d30, d31, d32, d33, e30, e31, e32, e33, f30, f31, f32, f33, g30, g31, g32, g33, h30, h31, h32, h33, i30, i31, i32, i33;
wire a40, a41, a42, a43, a44, a45, a46, a47, b40, b41, b42, b43, b44, b45, b46, b47, c40, c41, c42, c43, c44, c45, c46, c47, d40, d41, d42, d43, d44, d45, d46, d47, e40, e41, e42, e43, e44, e45, e46, e47, f40, f41, f42, f43, f44, f45, f46, f47, g40, g41, g42, g43, g44, g45, g46, g47, h40, h41, h42, h43, h44, h45, h46, h47, i40, i41, i42, i43, i44, i45, i46, i47;
wire m00, m01, m02, m03, m04, m05, m06, m07, m08, m09, m010, m011, m012, m013, m014, m015, n00, n01, n02, n03, n04, n05, n06, n07, n08, n09, n010, n011, n012, n013, n014, n015, o00, o01, o02, o03, o04, o05, o06, o07, o08, o09, o010, o011, o012, o013, o014, o015, p00, p01, p02, p03, p04, p05, p06, p07, p08, p09, p010, p011, p012, p013, p014, p015, q00, q01, q02, q03, q04, q05, q06, q07, q08, q09, q010, q011, q012, q013, q014, q015, r00, r01, r02, r03, r04, r05, r06, r07, r08, r09, r010, r011, r012, r013, r014, r015, s00, s01, s02, s03, s04, s05, s06, s07, s08, s09, s010, s011, s012, s013, s014, s015, t00, t01, t02, t03, t04, t05, t06, t07, t08, t09, t010, t011, t012, t013, t014, t015, u00, u01, u02, u03, u04, u05, u06, u07, u08, u09, u010, u011, u012, u013, u014, u015;
wire det0, det1, det2, det3, det4, det5, det6, det7, det8, det9, det10, det11, det12, det13, det14, det15, dummy;
wire as, bs, cs, ds, es, fs, gs, hs, is;

encoder1 encode1(a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, a23, a22, a21, a20);
encoder1 encode2(b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, b23, b22, b21, b20);
encoder1 encode3(c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, c23, c22, c21, c20);
encoder1 encode4(d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, d23, d22, d21, d20);
encoder1 encode5(e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, e23, e22, e21, e20);
encoder1 encode6(f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, f23, f22, f21, f20);
encoder1 encode7(g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, g23, g22, g21, g20);
encoder1 encode8(h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, h23, h22, h21, h20);
encoder1 encode9(i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, i23, i22, i21, i20);

encoder1 encode11(a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, a33, a32, a31, a30);
encoder1 encode12(b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, b33, b32, b31, b30);
encoder1 encode13(c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, c33, c32, c31, c30);
encoder1 encode14(d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, d33, d32, d31, d30);
encoder1 encode15(e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, e33, e32, e31, e30);
encoder1 encode16(f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, f33, f32, f31, f30);
encoder1 encode17(g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, g33, g32, g31, g30);
encoder1 encode18(h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, h33, h32, h31, h30);
encoder1 encode19(i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115, i33, i32, i31, i30);

det2 det21(e30, e31, e32, e33, f30, f31, f32, f33, h30, h31, h32, h33, i30, i31, i32, i33, a40, a41, a42, a43, a44, a45, a46, a47, as);
det2 det22(c30, c31, c32, c33, b30, b31, b32, b33, i30, i31, i32, i33, h30, h31, h32, h33, b40, b41, b42, b43, b44, b45, b46, b47, bs);
det2 det23(b30, b31, b32, b33, c30, c31, c32, c33, e30, e31, e32, e33, f30, f31, f32, f33, c40, c41, c42, c43, c44, c45, c46, c47, cs);
det2 det24(f30, f31, f32, f33, d30, d31, d32, d33, i30, i31, i32, i33, g30, g31, g32, g33, d40, d41, d42, d43, d44, d45, d46, d47, ds);
det2 det25(a30, a31, a32, a33, c30, c31, c32, c33, g30, g31, g32, g33, i30, i31, i32, i33, e40, e41, e42, e43, e44, e45, e46, e47, es);
det2 det26(c30, c31, c32, c33, a30, a31, a32, a33, f30, f31, f32, f33, d30, d31, d32, d33, f40, f41, f42, f43, f44, f45, f46, f47, fs);
det2 det27(d30, d31, d32, d33, e30, e31, e32, e33, g30, g31, g32, g33, h30, h31, h32, h33, g40, g41, g42, g43, g44, g45, g46, g47, gs);
det2 det28(b30, b31, b32, b33, a30, a31, a32, a33, h30, h31, h32, h33, g30, g31, g32, g33, h40, h41, h42, h43, h44, h45, h46, h47, hs);
det2 det29(a30, a31, a32, a33, b30, b31, b32, b33, d30, d31, d32, d33, e30, e31, e32, e33, i40, i41, i42, i43, i44, i45, i46, i47, is);

elements2 element1(a20, a21, a22, a23, b20, b21, b22, b23, c20, c21, c22, c23, a40, a41, a42, a43, a44, a45, a46, a47, as, d40, d41, d42, d43, d44, d45, d46, d47, ds, g40, g41, g42, g43, g44, g45, g46, g47, gs, m00, m01, m02, m03, m04, m05, m06, m07, m08, m09, m010, m011, m012, m013, m014, m015);
elements2 element2(a20, a21, a22, a23, b20, b21, b22, b23, c20, c21, c22, c23, b40, b41, b42, b43, b44, b45, b46, b47, bs, e40, e41, e42, e43, e44, e45, e46, e47, es, h40, h41, h42, h43, h44, h45, h46, h47, hs, n00, n01, n02, n03, n04, n05, n06, n07, n08, n09, n010, n011, n012, n013, n014, n015);
elements2 element3(a20, a21, a22, a23, b20, b21, b22, b23, c20, c21, c22, c23, c40, c41, c42, c43, c44, c45, c46, c47, cs, f40, f41, f42, f43, f44, f45, f46, f47, fs, i40, i41, i42, i43, i44, i45, i46, i47, is, o00, o01, o02, o03, o04, o05, o06, o07, o08, o09, o010, o011, o012, o013, o014, o015);
elements2 element4(d20, d21, d22, d23, e20, e21, e22, e23, f20, f21, f22, f23, a40, a41, a42, a43, a44, a45, a46, a47, as, d40, d41, d42, d43, d44, d45, d46, d47, ds, g40, g41, g42, g43, g44, g45, g46, g47, gs, p00, p01, p02, p03, p04, p05, p06, p07, p08, p09, p010, p011, p012, p013, p014, p015);
elements2 element5(d20, d21, d22, d23, e20, e21, e22, e23, f20, f21, f22, f23, b40, b41, b42, b43, b44, b45, b46, b47, bs, e40, e41, e42, e43, e44, e45, e46, e47, es, h40, h41, h42, h43, h44, h45, h46, h47, hs, q00, q01, q02, q03, q04, q05, q06, q07, q08, q09, q010, q011, q012, q013, q014, q015);
elements2 element6(d20, d21, d22, d23, e20, e21, e22, e23, f20, f21, f22, f23, c40, c41, c42, c43, c44, c45, c46, c47, cs, f40, f41, f42, f43, f44, f45, f46, f47, fs, i40, i41, i42, i43, i44, i45, i46, i47, is, r00, r01, r02, r03, r04, r05, r06, r07, r08, r09, r010, r011, r012, r013, r014, r015);
elements2 element7(g20, g21, g22, g23, h20, h21, h22, h33, i20, i21, i22, i23, a40, a41, a42, a43, a44, a45, a46, a47, as, d40, d41, d42, d43, d44, d45, d46, d47, ds, g40, g41, g42, g43, g44, g45, g46, g47, gs, s00, s01, s02, s03, s04, s05, s06, s07, s08, s09, s010, s011, s012, s013, s014, s015);
elements2 element8(g20, g21, g22, g23, h20, h21, h22, h23, i20, i21, i22, i23, b40, b41, b42, b43, b44, b45, b46, b47, bs, e40, e41, e42, e43, e44, e45, e46, e47, es, h40, h41, h42, h43, h44, h45, h46, h47, hs, t00, t01, t02, t03, t04, t05, t06, t07, t08, t09, t010, t011, t012, t013, t014, t015);
elements2 element9(g20, g21, g22, g23, h20, h21, h22, h23, i20, i21, i22, i23, c40, c41, c42, c43, c44, c45, c46, c47, cs, f40, f41, f42, f43, f44, f45, f46, f47, fs, i40, i41, i42, i43, i44, i45, i46, i47, is, u00, u01, u02, u03, u04, u05, u06, u07, u08, u09, u010, u011, u012, u013, u014, u015);

det3 det31(a30, a31, a32, a33, b30, b31, b32, b33, c30, c31, c32, c33, d30, d31, d32, d33, e30, e31, e32, e33, f30, f31, f32, f33, g30, g31, g32, g33, h30, h31, h32, h33, i30, i31, i32, i33, det0, det1, det2, det3, det4, det5, det6, det7, det8, det9, det10, det11, det12, det13, det14, det15);

division2 divide1(det0, det1, det2, det3, det4, det5, det6, det7, det8, det9, det10, det11, det12, det13, det14, 0, m00, m01, m02, m03, m04, m05, m06, m07, m08, m09, m010, m011, m012, m013, m014, m015, outa0, outa1, outa2, outa3, outa4, outa5, outa6, outa7, outa8, outa9, outa10, outa11, outa12, outa13, outa14, dummy);
division2 divide2(det0, det1, det2, det3, det4, det5, det6, det7, det8, det9, det10, det11, det12, det13, det14, 0, n00, n01, n02, n03, n04, n05, n06, n07, n08, n09, n010, n011, n012, n013, n014, n015, outb0, outb1, outb2, outb3, outb4, outb5, outb6, outb7, outb8, outb9, outb10, outb11, outb12, outb13, outb14, dummy);
division2 divide3(det0, det1, det2, det3, det4, det5, det6, det7, det8, det9, det10, det11, det12, det13, det14, 0, o00, o01, o02, o03, o04, o05, o06, o07, o08, o09, o010, o011, o012, o013, o014, o015, outc0, outc1, outc2, outc3, outc4, outc5, outc6, outc7, outc8, outc9, outc10, outc11, outc12, outc13, outc14, dummy);
division2 divide4(det0, det1, det2, det3, det4, det5, det6, det7, det8, det9, det10, det11, det12, det13, det14, 0, p00, p01, p02, p03, p04, p05, p06, p07, p08, p09, p010, p011, p012, p013, p014, p015, outd0, outd1, outd2, outd3, outd4, outd5, outd6, outd7, outd8, outd9, outd10, outd11, outd12, outd13, outd14, dummy);
division2 divide5(det0, det1, det2, det3, det4, det5, det6, det7, det8, det9, det10, det11, det12, det13, det14, 0, q00, q01, q02, q03, q04, q05, q06, q07, q08, q09, q010, q011, q012, q013, q014, q015, oute0, oute1, oute2, oute3, oute4, oute5, oute6, oute7, oute8, oute9, oute10, oute11, oute12, oute13, oute14, dummy);
division2 divide6(det0, det1, det2, det3, det4, det5, det6, det7, det8, det9, det10, det11, det12, det13, det14, 0, r00, r01, r02, r03, r04, r05, r06, r07, r08, r09, r010, r011, r012, r013, r014, r015, outf0, outf1, outf2, outf3, outf4, outf5, outf6, outf7, outf8, outf9, outf10, outf11, outf12, outf13, outf14, dummy);
division2 divide7(det0, det1, det2, det3, det4, det5, det6, det7, det8, det9, det10, det11, det12, det13, det14, 0, s00, s01, s02, s03, s04, s05, s06, s07, s08, s09, s010, s011, s012, s013, s014, s015, outg0, outg1, outg2, outg3, outg4, outg5, outg6, outg7, outg8, outg9, outg10, outg11, outg12, outg13, outg14, dummy);
division2 divide8(det0, det1, det2, det3, det4, det5, det6, det7, det8, det9, det10, det11, det12, det13, det14, 0, t00, t01, t02, t03, t04, t05, t06, t07, t08, t09, t010, t011, t012, t013, t014, t015, outh0, outh1, outh2, outh3, outh4, outh5, outh6, outh7, outh8, outh9, outh10, outh11, outh12, outh13, outh14, dummy);
division2 divide9(det0, det1, det2, det3, det4, det5, det6, det7, det8, det9, det10, det11, det12, det13, det14, 0, u00, u01, u02, u03, u04, u05, u06, u07, u08, u09, u010, u011, u012, u013, u014, u015, outi0, outi1, outi2, outi3, outi4, outi5, outi6, outi7, outi8, outi9, outi10, outi11, outi12, outi13, outi14, dummy);

or(outa15, det15, as);
or(outb15, det15, bs);
or(outc15, det15, cs);
or(outd15, det15, ds);
or(oute15, det15, es);
or(outf15, det15, fs);
or(outg15, det15, gs);
or(outh15, det15, hs);
or(outi15, det15, is);

endmodule
