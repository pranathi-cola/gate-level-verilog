module neo_matrix_tb;

reg choice2, choice1, choice0, a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115;
wire outa0, outa1, outa2, outa3, outa4, outa5, outa6, outa7, outa8, outa9, outa10, outa11, outa12, outa13, outa14, outa15, outb0, outb1, outb2, outb3, outb4, outb5, outb6, outb7, outb8, outb9, outb10, outb11, outb12, outb13, outb14, outb15, outc0, outc1, outc2, outc3, outc4, outc5, outc6, outc7, outc8, outc9, outc10, outc11, outc12, outc13, outc14, outc15, outd0, outd1, outd2, outd3, outd4, outd5, outd6, outd7, outd8, outd9, outd10, outd11, outd12, outd13, outd14, outd15, oute0, oute1, oute2, oute3, oute4, oute5, oute6, oute7, oute8, oute9, oute10, oute11, oute12, oute13, oute14, oute15, outf0, outf1, outf2, outf3, outf4, outf5, outf6, outf7, outf8, outf9, outf10, outf11, outf12, outf13, outf14, outf15, outg0, outg1, outg2, outg3, outg4, outg5, outg6, outg7, outg8, outg9, outg10, outg11, outg12, outg13, outg14, outg15, outh0, outh1, outh2, outh3, outh4, outh5, outh6, outh7, outh8, outh9, outh10, outh11, outh12, outh13, outh14, outh15, outi0, outi1, outi2, outi3, outi4, outi5, outi6, outi7, outi8, outi9, outi10, outi11, outi12, outi13, outi14, outi15;

neo_matrix matrixx1(choice2, choice1, choice0, a00, a01, a02, a03, a04, a05, a06, a07, a08, a09, a010, a011, a012, a013, a014, a015, b00, b01, b02, b03, b04, b05, b06, b07, b08, b09, b010, b011, b012, b013, b014, b015, c00, c01, c02, c03, c04, c05, c06, c07, c08, c09, c010, c011, c012, c013, c014, c015, d00, d01, d02, d03, d04, d05, d06, d07, d08, d09, d010, d011, d012, d013, d014, d015, e00, e01, e02, e03, e04, e05, e06, e07, e08, e09, e010, e011, e012, e013, e014, e015, f00, f01, f02, f03, f04, f05, f06, f07, f08, f09, f010, f011, f012, f013, f014, f015, g00, g01, g02, g03, g04, g05, g06, g07, g08, g09, g010, g011, g012, g013, g014, g015, h00, h01, h02, h03, h04, h05, h06, h07, h08, h09, h010, h011, h012, h013, h014, h015, i00, i01, i02, i03, i04, i05, i06, i07, i08, i09, i010, i011, i012, i013, i014, i015, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a110, a111, a112, a113, a114, a115, b10, b11, b12, b13, b14, b15, b16, b17, b18, b19, b110, b111, b112, b113, b114, b115, c10, c11, c12, c13, c14, c15, c16, c17, c18, c19, c110, c111, c112, c113, c114, c115, d10, d11, d12, d13, d14, d15, d16, d17, d18, d19, d110, d111, d112, d113, d114, d115, e10, e11, e12, e13, e14, e15, e16, e17, e18, e19, e110, e111, e112, e113, e114, e115, f10, f11, f12, f13, f14, f15, f16, f17, f18, f19, f110, f111, f112, f113, f114, f115, g10, g11, g12, g13, g14, g15, g16, g17, g18, g19, g110, g111, g112, g113, g114, g115, h10, h11, h12, h13, h14, h15, h16, h17, h18, h19, h110, h111, h112, h113, h114, h115, i10, i11, i12, i13, i14, i15, i16, i17, i18, i19, i110, i111, i112, i113, i114, i115, outa0, outa1, outa2, outa3, outa4, outa5, outa6, outa7, outa8, outa9, outa10, outa11, outa12, outa13, outa14, outa15, outb0, outb1, outb2, outb3, outb4, outb5, outb6, outb7, outb8, outb9, outb10, outb11, outb12, outb13, outb14, outb15, outc0, outc1, outc2, outc3, outc4, outc5, outc6, outc7, outc8, outc9, outc10, outc11, outc12, outc13, outc14, outc15, outd0, outd1, outd2, outd3, outd4, outd5, outd6, outd7, outd8, outd9, outd10, outd11, outd12, outd13, outd14, outd15, oute0, oute1, oute2, oute3, oute4, oute5, oute6, oute7, oute8, oute9, oute10, oute11, oute12, oute13, oute14, oute15, outf0, outf1, outf2, outf3, outf4, outf5, outf6, outf7, outf8, outf9, outf10, outf11, outf12, outf13, outf14, outf15, outg0, outg1, outg2, outg3, outg4, outg5, outg6, outg7, outg8, outg9, outg10, outg11, outg12, outg13, outg14, outg15, outh0, outh1, outh2, outh3, outh4, outh5, outh6, outh7, outh8, outh9, outh10, outh11, outh12, outh13, outh14, outh15, outi0, outi1, outi2, outi3, outi4, outi5, outi6, outi7, outi8, outi9, outi10, outi11, outi12, outi13, outi14, outi15);

initial begin

#5
choice2=0; choice1=0; choice0=0; a00=0; a01=0; a02=0; a03=0; a04=0; a05=0; a06=0; a07=1; a08=0; a09=0; a010=0; a011=0; a012=0; a013=0; a014=0; a015=0; b00=0; b01=0; b02=0; b03=0; b04=1; b05=0; b06=0; b07=0; b08=0; b09=0; b010=0; b011=0; b012=0; b013=0; b014=0; b015=0; c00=0; c01=0; c02=0; c03=0; c04=0; c05=0; c06=0; c07=1; c08=0; c09=0; c010=0; c011=0; c012=0; c013=0; c014=0; c015=0; d00=0; d01=0; d02=0; d03=1; d04=0; d05=0; d06=0; d07=0; d08=0; d09=0; d010=0; d011=0; d012=0; d013=0; d014=0; d015=0; e00=0; e01=1; e02=0; e03=0; e04=0; e05=0; e06=0; e07=0; e08=0; e09=0; e010=0; e011=0; e012=0; e013=0; e014=0; e015=0; f00=1; f01=0; f02=0; f03=0; f04=0; f05=0; f06=0; f07=0; f08=0; f09=0; f010=0; f011=0; f012=0; f013=0; f014=0; f015=0; g00=0; g01=1; g02=0; g03=0; g04=0; g05=0; g06=0; g07=0; g08=0; g09=0; g010=0; g011=0; g012=0; g013=0; g014=0; g015=0; h00=0; h01=0; h02=0; h03=0; h04=1; h05=0; h06=0; h07=0; h08=0; h09=0; h010=0; h011=0; h012=0; h013=0; h014=0; h015=0; i00=0; i01=1; i02=0; i03=0; i04=0; i05=0; i06=0; i07=0; i08=0; i09=0; i010=0; i011=0; i012=0; i013=0; i014=0; i015=0; a10=0; a11=0; a12=1; a13=0; a14=0; a15=0; a16=0; a17=0; a18=0; a19=0; a110=0; a111=0; a112=0; a113=0; a114=0; a115=0; b10=0; b11=1; b12=0; b13=0; b14=0; b15=0; b16=0; b17=0; b18=0; b19=0; b110=0; b111=0; b112=0; b113=0; b114=0; b115=0; c10=1; c11=0; c12=0; c13=0; c14=0; c15=0; c16=0; c17=0; c18=0; c19=0; c110=0; c111=0; c112=0; c113=0; c114=0; c115=0; d10=1; d11=0; d12=0; d13=0; d14=0; d15=0; d16=0; d17=0; d18=0; d19=0; d110=0; d111=0; d112=0; d113=0; d114=0; d115=0; e10=1; e11=0; e12=0; e13=0; e14=0; e15=0; e16=0; e17=0; e18=0; e19=0; e110=0; e111=0; e112=0; e113=0; e114=0; e115=0; f10=1; f11=0; f12=0; f13=0; f14=0; f15=0; f16=0; f17=0; f18=0; f19=0; f110=0; f111=0; f112=0; f113=0; f114=0; f115=0; g10=0; g11=0; g12=1; g13=0; g14=0; g15=0; g16=0; g17=0; g18=0; g19=0; g110=0; g111=0; g112=0; g113=0; g114=0; g115=0; h10=0; h11=0; h12=0; h13=0; h14=0; h15=0; h16=0; h17=0; h18=0; h19=1; h110=0; h111=0; h112=0; h113=0; h114=0; h115=0; i10=0; i11=1; i12=0; i13=0; i14=0; i15=0; i16=0; i17=0; i18=0; i19=0; i110=0; i111=0; i112=0; i113=0; i114=0; i115=0;
#500
choice2=0; choice1=0; choice0=1; a00=0; a01=0; a02=0; a03=0; a04=0; a05=0; a06=0; a07=1; a08=0; a09=0; a010=0; a011=0; a012=0; a013=0; a014=0; a015=0; b00=0; b01=0; b02=0; b03=0; b04=1; b05=0; b06=0; b07=0; b08=0; b09=0; b010=0; b011=0; b012=0; b013=0; b014=0; b015=0; c00=0; c01=0; c02=0; c03=0; c04=0; c05=0; c06=0; c07=1; c08=0; c09=0; c010=0; c011=0; c012=0; c013=0; c014=0; c015=0; d00=0; d01=0; d02=0; d03=1; d04=0; d05=0; d06=0; d07=0; d08=0; d09=0; d010=0; d011=0; d012=0; d013=0; d014=0; d015=0; e00=0; e01=1; e02=0; e03=0; e04=0; e05=0; e06=0; e07=0; e08=0; e09=0; e010=0; e011=0; e012=0; e013=0; e014=0; e015=0; f00=1; f01=0; f02=0; f03=0; f04=0; f05=0; f06=0; f07=0; f08=0; f09=0; f010=0; f011=0; f012=0; f013=0; f014=0; f015=0; g00=0; g01=1; g02=0; g03=0; g04=0; g05=0; g06=0; g07=0; g08=0; g09=0; g010=0; g011=0; g012=0; g013=0; g014=0; g015=0; h00=0; h01=0; h02=0; h03=0; h04=1; h05=0; h06=0; h07=0; h08=0; h09=0; h010=0; h011=0; h012=0; h013=0; h014=0; h015=0; i00=0; i01=1; i02=0; i03=0; i04=0; i05=0; i06=0; i07=0; i08=0; i09=0; i010=0; i011=0; i012=0; i013=0; i014=0; i015=0; a10=0; a11=0; a12=1; a13=0; a14=0; a15=0; a16=0; a17=0; a18=0; a19=0; a110=0; a111=0; a112=0; a113=0; a114=0; a115=0; b10=0; b11=1; b12=0; b13=0; b14=0; b15=0; b16=0; b17=0; b18=0; b19=0; b110=0; b111=0; b112=0; b113=0; b114=0; b115=0; c10=1; c11=0; c12=0; c13=0; c14=0; c15=0; c16=0; c17=0; c18=0; c19=0; c110=0; c111=0; c112=0; c113=0; c114=0; c115=0; d10=1; d11=0; d12=0; d13=0; d14=0; d15=0; d16=0; d17=0; d18=0; d19=0; d110=0; d111=0; d112=0; d113=0; d114=0; d115=0; e10=1; e11=0; e12=0; e13=0; e14=0; e15=0; e16=0; e17=0; e18=0; e19=0; e110=0; e111=0; e112=0; e113=0; e114=0; e115=0; f10=1; f11=0; f12=0; f13=0; f14=0; f15=0; f16=0; f17=0; f18=0; f19=0; f110=0; f111=0; f112=0; f113=0; f114=0; f115=0; g10=0; g11=0; g12=1; g13=0; g14=0; g15=0; g16=0; g17=0; g18=0; g19=0; g110=0; g111=0; g112=0; g113=0; g114=0; g115=0; h10=0; h11=0; h12=0; h13=0; h14=0; h15=0; h16=0; h17=0; h18=0; h19=1; h110=0; h111=0; h112=0; h113=0; h114=0; h115=0; i10=0; i11=1; i12=0; i13=0; i14=0; i15=0; i16=0; i17=0; i18=0; i19=0; i110=0; i111=0; i112=0; i113=0; i114=0; i115=0;
#500
choice2=0; choice1=1; choice0=0; a00=0; a01=0; a02=0; a03=0; a04=0; a05=0; a06=0; a07=1; a08=0; a09=0; a010=0; a011=0; a012=0; a013=0; a014=0; a015=0; b00=0; b01=0; b02=0; b03=0; b04=1; b05=0; b06=0; b07=0; b08=0; b09=0; b010=0; b011=0; b012=0; b013=0; b014=0; b015=0; c00=0; c01=0; c02=0; c03=0; c04=0; c05=0; c06=0; c07=1; c08=0; c09=0; c010=0; c011=0; c012=0; c013=0; c014=0; c015=0; d00=0; d01=0; d02=0; d03=1; d04=0; d05=0; d06=0; d07=0; d08=0; d09=0; d010=0; d011=0; d012=0; d013=0; d014=0; d015=0; e00=0; e01=1; e02=0; e03=0; e04=0; e05=0; e06=0; e07=0; e08=0; e09=0; e010=0; e011=0; e012=0; e013=0; e014=0; e015=0; f00=1; f01=0; f02=0; f03=0; f04=0; f05=0; f06=0; f07=0; f08=0; f09=0; f010=0; f011=0; f012=0; f013=0; f014=0; f015=0; g00=0; g01=1; g02=0; g03=0; g04=0; g05=0; g06=0; g07=0; g08=0; g09=0; g010=0; g011=0; g012=0; g013=0; g014=0; g015=0; h00=0; h01=0; h02=0; h03=0; h04=1; h05=0; h06=0; h07=0; h08=0; h09=0; h010=0; h011=0; h012=0; h013=0; h014=0; h015=0; i00=0; i01=1; i02=0; i03=0; i04=0; i05=0; i06=0; i07=0; i08=0; i09=0; i010=0; i011=0; i012=0; i013=0; i014=0; i015=0; a10=0; a11=0; a12=1; a13=0; a14=0; a15=0; a16=0; a17=0; a18=0; a19=0; a110=0; a111=0; a112=0; a113=0; a114=0; a115=0; b10=0; b11=1; b12=0; b13=0; b14=0; b15=0; b16=0; b17=0; b18=0; b19=0; b110=0; b111=0; b112=0; b113=0; b114=0; b115=0; c10=1; c11=0; c12=0; c13=0; c14=0; c15=0; c16=0; c17=0; c18=0; c19=0; c110=0; c111=0; c112=0; c113=0; c114=0; c115=0; d10=1; d11=0; d12=0; d13=0; d14=0; d15=0; d16=0; d17=0; d18=0; d19=0; d110=0; d111=0; d112=0; d113=0; d114=0; d115=0; e10=1; e11=0; e12=0; e13=0; e14=0; e15=0; e16=0; e17=0; e18=0; e19=0; e110=0; e111=0; e112=0; e113=0; e114=0; e115=0; f10=1; f11=0; f12=0; f13=0; f14=0; f15=0; f16=0; f17=0; f18=0; f19=0; f110=0; f111=0; f112=0; f113=0; f114=0; f115=0; g10=0; g11=0; g12=1; g13=0; g14=0; g15=0; g16=0; g17=0; g18=0; g19=0; g110=0; g111=0; g112=0; g113=0; g114=0; g115=0; h10=0; h11=0; h12=0; h13=0; h14=0; h15=0; h16=0; h17=0; h18=0; h19=1; h110=0; h111=0; h112=0; h113=0; h114=0; h115=0; i10=0; i11=1; i12=0; i13=0; i14=0; i15=0; i16=0; i17=0; i18=0; i19=0; i110=0; i111=0; i112=0; i113=0; i114=0; i115=0;
#500
choice2=0; choice1=1; choice0=1; a00=0; a01=0; a02=0; a03=0; a04=0; a05=0; a06=0; a07=1; a08=0; a09=0; a010=0; a011=0; a012=0; a013=0; a014=0; a015=0; b00=0; b01=0; b02=0; b03=0; b04=1; b05=0; b06=0; b07=0; b08=0; b09=0; b010=0; b011=0; b012=0; b013=0; b014=0; b015=0; c00=0; c01=0; c02=0; c03=0; c04=0; c05=0; c06=0; c07=1; c08=0; c09=0; c010=0; c011=0; c012=0; c013=0; c014=0; c015=0; d00=0; d01=0; d02=0; d03=1; d04=0; d05=0; d06=0; d07=0; d08=0; d09=0; d010=0; d011=0; d012=0; d013=0; d014=0; d015=0; e00=0; e01=1; e02=0; e03=0; e04=0; e05=0; e06=0; e07=0; e08=0; e09=0; e010=0; e011=0; e012=0; e013=0; e014=0; e015=0; f00=1; f01=0; f02=0; f03=0; f04=0; f05=0; f06=0; f07=0; f08=0; f09=0; f010=0; f011=0; f012=0; f013=0; f014=0; f015=0; g00=0; g01=1; g02=0; g03=0; g04=0; g05=0; g06=0; g07=0; g08=0; g09=0; g010=0; g011=0; g012=0; g013=0; g014=0; g015=0; h00=0; h01=0; h02=0; h03=0; h04=1; h05=0; h06=0; h07=0; h08=0; h09=0; h010=0; h011=0; h012=0; h013=0; h014=0; h015=0; i00=0; i01=1; i02=0; i03=0; i04=0; i05=0; i06=0; i07=0; i08=0; i09=0; i010=0; i011=0; i012=0; i013=0; i014=0; i015=0; a10=0; a11=0; a12=1; a13=0; a14=0; a15=0; a16=0; a17=0; a18=0; a19=0; a110=0; a111=0; a112=0; a113=0; a114=0; a115=0; b10=0; b11=1; b12=0; b13=0; b14=0; b15=0; b16=0; b17=0; b18=0; b19=0; b110=0; b111=0; b112=0; b113=0; b114=0; b115=0; c10=1; c11=0; c12=0; c13=0; c14=0; c15=0; c16=0; c17=0; c18=0; c19=0; c110=0; c111=0; c112=0; c113=0; c114=0; c115=0; d10=1; d11=0; d12=0; d13=0; d14=0; d15=0; d16=0; d17=0; d18=0; d19=0; d110=0; d111=0; d112=0; d113=0; d114=0; d115=0; e10=1; e11=0; e12=0; e13=0; e14=0; e15=0; e16=0; e17=0; e18=0; e19=0; e110=0; e111=0; e112=0; e113=0; e114=0; e115=0; f10=1; f11=0; f12=0; f13=0; f14=0; f15=0; f16=0; f17=0; f18=0; f19=0; f110=0; f111=0; f112=0; f113=0; f114=0; f115=0; g10=0; g11=0; g12=1; g13=0; g14=0; g15=0; g16=0; g17=0; g18=0; g19=0; g110=0; g111=0; g112=0; g113=0; g114=0; g115=0; h10=0; h11=0; h12=0; h13=0; h14=0; h15=0; h16=0; h17=0; h18=0; h19=1; h110=0; h111=0; h112=0; h113=0; h114=0; h115=0; i10=0; i11=1; i12=0; i13=0; i14=0; i15=0; i16=0; i17=0; i18=0; i19=0; i110=0; i111=0; i112=0; i113=0; i114=0; i115=0;
#500
choice2=1; choice1=0; choice0=0; a00=0; a01=0; a02=0; a03=0; a04=0; a05=0; a06=0; a07=1; a08=0; a09=0; a010=0; a011=0; a012=0; a013=0; a014=0; a015=0; b00=0; b01=0; b02=0; b03=0; b04=1; b05=0; b06=0; b07=0; b08=0; b09=0; b010=0; b011=0; b012=0; b013=0; b014=0; b015=0; c00=0; c01=0; c02=0; c03=0; c04=0; c05=0; c06=0; c07=1; c08=0; c09=0; c010=0; c011=0; c012=0; c013=0; c014=0; c015=0; d00=0; d01=0; d02=0; d03=1; d04=0; d05=0; d06=0; d07=0; d08=0; d09=0; d010=0; d011=0; d012=0; d013=0; d014=0; d015=0; e00=0; e01=1; e02=0; e03=0; e04=0; e05=0; e06=0; e07=0; e08=0; e09=0; e010=0; e011=0; e012=0; e013=0; e014=0; e015=0; f00=1; f01=0; f02=0; f03=0; f04=0; f05=0; f06=0; f07=0; f08=0; f09=0; f010=0; f011=0; f012=0; f013=0; f014=0; f015=0; g00=0; g01=1; g02=0; g03=0; g04=0; g05=0; g06=0; g07=0; g08=0; g09=0; g010=0; g011=0; g012=0; g013=0; g014=0; g015=0; h00=0; h01=0; h02=0; h03=0; h04=1; h05=0; h06=0; h07=0; h08=0; h09=0; h010=0; h011=0; h012=0; h013=0; h014=0; h015=0; i00=0; i01=1; i02=0; i03=0; i04=0; i05=0; i06=0; i07=0; i08=0; i09=0; i010=0; i011=0; i012=0; i013=0; i014=0; i015=0; a10=0; a11=0; a12=1; a13=0; a14=0; a15=0; a16=0; a17=0; a18=0; a19=0; a110=0; a111=0; a112=0; a113=0; a114=0; a115=0; b10=0; b11=1; b12=0; b13=0; b14=0; b15=0; b16=0; b17=0; b18=0; b19=0; b110=0; b111=0; b112=0; b113=0; b114=0; b115=0; c10=1; c11=0; c12=0; c13=0; c14=0; c15=0; c16=0; c17=0; c18=0; c19=0; c110=0; c111=0; c112=0; c113=0; c114=0; c115=0; d10=1; d11=0; d12=0; d13=0; d14=0; d15=0; d16=0; d17=0; d18=0; d19=0; d110=0; d111=0; d112=0; d113=0; d114=0; d115=0; e10=1; e11=0; e12=0; e13=0; e14=0; e15=0; e16=0; e17=0; e18=0; e19=0; e110=0; e111=0; e112=0; e113=0; e114=0; e115=0; f10=1; f11=0; f12=0; f13=0; f14=0; f15=0; f16=0; f17=0; f18=0; f19=0; f110=0; f111=0; f112=0; f113=0; f114=0; f115=0; g10=0; g11=0; g12=1; g13=0; g14=0; g15=0; g16=0; g17=0; g18=0; g19=0; g110=0; g111=0; g112=0; g113=0; g114=0; g115=0; h10=0; h11=0; h12=0; h13=0; h14=0; h15=0; h16=0; h17=0; h18=0; h19=1; h110=0; h111=0; h112=0; h113=0; h114=0; h115=0; i10=0; i11=1; i12=0; i13=0; i14=0; i15=0; i16=0; i17=0; i18=0; i19=0; i110=0; i111=0; i112=0; i113=0; i114=0; i115=0;
#500;

end 

endmodule
